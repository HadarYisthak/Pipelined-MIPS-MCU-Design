---------------------------------------------------------------------------------------------
-- Copyright 2025 Hananya Ribo 
-- Advanced CPU architecture and Hardware Accelerators Lab 361-1-4693 BGU
---------------------------------------------------------------------------------------------
--  Idecode module (implements the register file for the MIPS computer
LIBRARY IEEE; 		
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY Idecode IS
	generic(
		DATA_BUS_WIDTH : integer := 32
	);
	PORT(		clk_i,rst_i			: IN 	STD_LOGIC;
			instruction_i 			: IN 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			RegWrite_ctrl_i 		: IN 	STD_LOGIC;
			Jump				: IN	STD_LOGIC;
			pc_plus_4_i			: IN	STD_LOGIC_VECTOR(7 DOWNTO 0);
			ForwardA_ID, ForwardB_ID	: IN 	STD_LOGIC;
			write_register_address      	: IN    STD_LOGIC_VECTOR(4 DOWNTO 0);
			Branch_read_data_FW		: IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
			Branch_ctrl_i			: IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
			Stall_ID			: IN    STD_LOGIC;
			write_reg_data_i		: IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
			PCSrc		 		: OUT 	STD_LOGIC_VECTOR(1 DOWNTO 0);
			read_data_1_o			: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			read_data_2_o			: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			sign_extend_o 			: OUT 	STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
			read_register_1_address_w 	: OUT 	STD_LOGIC_VECTOR(4 DOWNTO 0);
			read_register_2_address_w 	: OUT 	STD_LOGIC_VECTOR(4 DOWNTO 0);
			write_register_address_0 	: OUT 	STD_LOGIC_VECTOR(4 DOWNTO 0);
			write_register_address_1 	: OUT 	STD_LOGIC_VECTOR(4 DOWNTO 0);
			pc_jump_o			: OUT   STD_LOGIC_VECTOR(7 DOWNTO 0);
			pc_branch_o 			: OUT 	STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END Idecode;


ARCHITECTURE behavior OF Idecode IS
TYPE register_file IS ARRAY (0 TO 31) OF STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);

	SIGNAL RF_q				: register_file;
	SIGNAL rd_register_w, read_register_1_address_sig, read_register_2_address_sig: STD_LOGIC_VECTOR( 4 DOWNTO 0 );
	SIGNAL imm_value_w			: STD_LOGIC_VECTOR( 15 DOWNTO 0 );
	SIGNAL read_data_1_sig, read_data_2_sig	: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL comp_1_w, comp_2_w		: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL Sign_extend_sig 			: STD_LOGIC_VECTOR( 31 DOWNTO 0 );

BEGIN
-------????? ???? ???????
	read_register_1_address_w 	<= instruction_i(25 DOWNTO 21);
   	read_register_2_address_w 	<= instruction_i(20 DOWNTO 16);
	write_register_address_0 	<= Instruction_i(20 DOWNTO 16);
   	write_register_address_1	<= instruction_i(15 DOWNTO 11);
   	imm_value_w 			<= instruction_i(15 DOWNTO 0);
		read_register_1_address_sig <= read_register_1_address_w;
		read_register_2_address_sig <= read_register_2_address_w;

	-------------- Read Register 1 Operation ---------------------------
	comp_1_w  		<= read_data_1_sig WHEN ForwardA_ID = '0' ELSE Branch_read_data_FW;
	read_data_1_sig		<= RF_q(CONV_INTEGER(read_register_1_address_sig));
	read_data_1_o 		<= read_data_1_sig;
	-------------- Read Register 2 Operation ---------------------------		 
	comp_2_w 		<= read_data_2_sig WHEN ForwardB_ID = '0' ELSE Branch_read_data_FW;
	read_data_2_sig 	<= RF_q(CONV_INTEGER(read_register_2_address_sig));
	read_data_2_o 		<= read_data_2_sig;

	-------------- PCSrc from Read Register Comp -----------------------
	PCSrc(1) 		<= Jump;
	PCSrc(0) 		<= Branch_ctrl_i(0) WHEN ((comp_1_w = comp_2_w) AND Stall_ID = '0') ELSE 
				   Branch_ctrl_i(1) WHEN ((comp_1_w /= comp_2_w) AND Stall_ID = '0') ELSE '0';  -- Branch Comperator (For bne chen inequality)
	

		-------------  Calc PC Address when branching --------------------
	pc_branch_o 	<= 	pc_plus_4_i +  Sign_extend_sig(7 DOWNTO 0);
	pc_jump_o	<= 	Sign_extend_sig(7 DOWNTO 0) WHEN instruction_i(27) = '1' ELSE
				read_data_1_sig(7 DOWNTO 0); -- jr

	-------------- Sign Extend 16-bits to 32-bits ----------------------
    	Sign_extend_sig <= 	X"0000" & imm_value_w WHEN imm_value_w(15) = '0' ELSE
				X"FFFF" & imm_value_w;
	Sign_extend_o 	<=	Sign_extend_sig;

	----------- Register File Process ---------------
	process(clk_i,rst_i)
	begin
		if (rst_i='1') then
			FOR i IN 0 TO 31 LOOP
				-- RF_q(i) <= CONV_STD_LOGIC_VECTOR(i,32);
				RF_q(i) <= CONV_STD_LOGIC_VECTOR(0,32);
			END LOOP;
		elsif (clk_i'event and clk_i='0') then --write to RF in falling edge
			if (RegWrite_ctrl_i = '1' AND CONV_INTEGER(write_register_address) /= 0) then
				RF_q(CONV_INTEGER(CONV_INTEGER(write_register_address))) <= write_reg_data_i;
				-- index is integer type so we must use conv_integer for type casting
			end if;
		end if;
end process;

END behavior;





