library IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
use ieee.std_logic_unsigned.all;
USE work.aux_package.all;


ENTITY  ALU IS
	generic(
		DATA_BUS_WIDTH : integer := 32
	);
	PORT(		a_input_w 			: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			b_input_w 			: IN 	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
			ALU_ctl		 		: IN 	STD_LOGIC_VECTOR( 3 DOWNTO 0 );
			zero_o 				: OUT	STD_LOGIC;
			alu_res_o			: OUT   STD_LOGIC_VECTOR( 31 DOWNTO 0 )
			);
END ALU;
------------ Architecture -----------------
ARCHITECTURE behavior OF ALU IS

SIGNAL alu_out_mux_w		: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
SIGNAL shift_res_w		: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);
SIGNAL dir_w			:STD_LOGIC;
SIGNAL b_input_b		: STD_LOGIC_VECTOR(DATA_BUS_WIDTH-1 DOWNTO 0);

BEGIN
-- Generate Zero Flag
	zero_o <= 	'1' WHEN (alu_out_mux_w(DATA_BUS_WIDTH-1 DOWNTO 0) = X"00000000") ELSE
			'0'; 

-- Select ALU output        
	alu_res_o <= 	X"0000000" & B"000"  & alu_out_mux_w(31) WHEN  ALU_ctl = "0111" ELSE 
					alu_out_mux_w(DATA_BUS_WIDTH-1 DOWNTO 0);



---shifter---
dir_w 	<= 	'1' when ALU_ctl = "0101" ELSE
		'0';

b_input_b <=	(others => '0') WHEN (not(ALU_ctl="0101" or ALU_ctl="1000")) ELSE
		b_input_w;

shift_action : Shifter 
	GENERIC MAP(n=>  DATA_BUS_WIDTH)
	PORT MAP (
		y	=>	a_input_w,
		x	=>	b_input_b,
		dir	=>	dir_w,
		res	=>	shift_res_w
		);

PROCESS ( ALU_ctl, a_input_w, b_input_w )
	variable product : STD_LOGIC_VECTOR(63 downto 0); 
	BEGIN
	--------------- Select ALU operation ---------------------
 	CASE ALU_ctl IS
		-- ALU performs ALUresult = A_input AND B_input
		WHEN "0000" 	=>	alu_out_mux_w	<= a_input_w AND b_input_w ; 
		-- ALU performs ALUresult = A_input OR B_input
     		WHEN "0001" 	=>	alu_out_mux_w	<= a_input_w OR b_input_w ;
		-- ALU performs ALUresult = A_input + B_input
	 	WHEN "0010" 	=>	alu_out_mux_w 	<= a_input_w + b_input_w ; 
		-- ALU performs ALUresult = A_input * B_input
 	 	WHEN "0011" 	=>	product := a_input_w * b_input_w ; -- result 64 bit
							alu_out_mux_w <= product(31 DOWNTO 0); -- Take Lower Part
		-- ALU performs ALUresult = A_input XOR B_input
 	 	WHEN "0100" 	=>	alu_out_mux_w 	<= a_input_w XOR b_input_w ;
		-- ALU performs ALUresult = A_input SLL B_input
 	 	WHEN "0101" 	=>	alu_out_mux_w 	<=	shift_res_w;

		-- ALU performs ALUresult = A_input SRL B_input
 	 	WHEN "1000" 	=>	alu_out_mux_w 	<=	shift_res_w; 

		-- ALU performs ALUresult = A_input -B_input
 	 	WHEN "0110" 	=>	alu_out_mux_w 	<= a_input_w - b_input_w ; 
		-- ALU performs SLT
  	 	WHEN "0111" 	=>	alu_out_mux_w 	<= a_input_w - b_input_w ;  
		-- ALU performs LUI
  	 	WHEN "1001" 	=>	alu_out_mux_w 	<= b_input_w (15 DOWNTO 0) & "0000000000000000";
		-- ALU performs ADDU
  	 	WHEN "1101"	=>	alu_out_mux_w <= conv_std_logic_vector(unsigned(a_input_w) + unsigned(b_input_w), DATA_BUS_WIDTH);

		-- OUTPUT ZERO
 	 	WHEN OTHERS	=>	alu_out_mux_w 	<= X"00000000" ;
  	END CASE;
  END PROCESS;
END behavior;